** Generated for: hspiceD
** Generated on: Feb 19 15:12:42 2019
** Design library name: ET710_ADC_bhv
** Design cell name: TOP_IADC_1b_bhv
** Design view name: schematic


** Library name: ET710_ADC_bhv
** Cell name: fdopb
** View name: schematic
*.subckt fdopb agnd avdd inn inp ir on op pdn vcm vcmfb
*.ends fdopb
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: TGB
** View name: schematic
*.subckt TGB bi1 bi2 pwra sub t tn
*.ends TGB
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: dac_int_1bit
** View name: schematic
.subckt dac_int_1bit agnd avdd dacn dacp pvrefn pvrefn_b pvrefp pvrefp_b vrefn vrefp
xi6 vrefn dacn avdd agnd pvrefp pvrefp_b TGB
xi7 vrefp dacn avdd agnd pvrefn pvrefn_b TGB
xi40 vrefp dacp avdd agnd pvrefp pvrefp_b TGB
xi41 vrefn dacp avdd agnd pvrefn pvrefn_b TGB
.ends dac_int_1bit
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: int1_1b_bhv
** View name: schematic
.subckt int1_1b_bhv agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b inn inp iref outn outp pdn pvrefn pvrefn_b pvrefp pvrefp_b rst rst_b vcm vrefn vrefp
xop agnd avdd opin opip iref outn outp pdn vcm vcm fdopb
xdac agnd avdd dacn dacp pvrefn pvrefn_b pvrefp pvrefp_b vrefn vrefp dac_int_1bit
xswinn_0 inn dacn avdd agnd p1d p1d_b TGB
xswinn_1 inn dacn avdd agnd p1d p1d_b TGB
xswinn_2 inn dacn avdd agnd p1d p1d_b TGB
xswinn_3 inn dacn avdd agnd p1d p1d_b TGB
xswrst2 opip outn avdd agnd rst rst_b TGB
xsw6 cinn opip avdd agnd p2 p2_b TGB
xswrst1 opin outp avdd agnd rst rst_b TGB
xsw2 cinp opin avdd agnd p2 p2_b TGB
xsw3 vcm cinp avdd agnd p1 p1_b TGB
xswinp_0 inp dacp avdd agnd p1d p1d_b TGB
xswinp_1 inp dacp avdd agnd p1d p1d_b TGB
xswinp_2 inp dacp avdd agnd p1d p1d_b TGB
xswinp_3 inp dacp avdd agnd p1d p1d_b TGB
xsw7 vcm cinn avdd agnd p1 p1_b TGB
cfbp_1 opin outp 20e-15
cfbp_2 opin outp 20e-15
cfbp_3 opin outp 20e-15
cfbn_1 opip outn 20e-15
cfbn_2 opip outn 20e-15
cfbn_3 opip outn 20e-15
csn cinn dacn 20e-15
csp cinp dacp 20e-15
.ends int1_1b_bhv
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: PMOS_B
** View name: schematic
*.subckt PMOS_B b d g s
*.ends PMOS_B
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: NMOS_B
** View name: schematic
*.subckt NMOS_B b d g s
*.ends NMOS_B
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: inv_bhv
** View name: schematic
.subckt inv_bhv dgnd vdd y yn
r1 net23 yn 10
c1 yn dgnd 5e-15
xp1 vdd net23 y vdd PMOS_B
xn1 dgnd net23 y dgnd NMOS_B
.ends inv_bhv
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: nand2_bhv
** View name: schematic
.subckt nand2_bhv dgnd vdd y1 y2 yn
xn1 dgnd yn y2 net8 NMOS_B
xi9 dgnd net8 y1 dgnd NMOS_B
xp1 vdd yn y1 vdd PMOS_B
xi10 vdd yn y2 vdd PMOS_B
.ends nand2_bhv
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: clk_fb_1bit
** View name: schematic
.subckt clk_fb_1bit agnd avdd d p2 pvrefn pvrefn_b pvrefp pvrefp_b
xi64 agnd avdd pvrefn pvrefn_b inv_bhv
xi20 agnd avdd net43 pvrefp inv_bhv
xi60 agnd avdd net48 pvrefn inv_bhv
xi59 agnd avdd d d_b inv_bhv
xi63 agnd avdd pvrefp pvrefp_b inv_bhv
xi62 agnd avdd p2 d_b net48 nand2_bhv
xi19 agnd avdd p2 d net43 nand2_bhv
.ends clk_fb_1bit
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: preamp_cmp_b
** View name: schematic
*.subckt preamp_cmp_b agnd avdd inn inp ir on op pdn vcm vcmfb
*.ends preamp_cmp_b
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: Dlatch
** View name: schematic
.subckt Dlatch q d clk clkb dvdd dgnd
xi2 dgnd dvdd net017 q inv_bhv
xi1 dgnd dvdd net22 net8 inv_bhv
c0 q dgnd 5e-15
c1 net017 dgnd 5e-15
r1 net8 net017 2
xi29 d net22 dvdd dgnd clk clkb TGB
xsw1 net22 q dvdd dgnd clkb clk TGB
.ends Dlatch
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: dff
** View name: schematic
.subckt dff q d clk clkb dvdd dgnd
xi13 net275 d clkb clk dvdd dgnd Dlatch
xi14 q net275 clk clkb dvdd dgnd Dlatch
.ends dff
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: amp_cmp
** View name: schematic
*.subckt amp_cmp vm vout vp
*.ends amp_cmp
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: cmp_clk
** View name: schematic
.subckt cmp_clk agnd avdd clk clk_b inn inp y
xdff y net22 clk clk_b avdd agnd dff
xpreamp inn net22 inp amp_cmp
.ends cmp_clk
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: adder_cmp_1b_CIFF2
** View name: schematic
.subckt adder_cmp_1b_CIFF2 agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b d iref pdn uin_n uin_p vcm vthn vthp int1n int1p int2n int2p
xpreamp_bhv agnd avdd opin opip iref amp_n amp_p pdn vcm vcm preamp_cmp_b
xcmp3 agnd avdd p1_b p1 amp_n amp_p d_b cmp_clk
xi1 agnd avdd d_b d inv_bhv
xi52 amp_p opin avdd agnd p2 p2_b TGB
xi63 vcm net088 avdd agnd p2d p2d_b TGB
xi62 uin_p net088 avdd agnd p1d p1d_b TGB
xi55 int1p net0107 avdd agnd p1d p1d_b TGB
xi56 vcm net0107 avdd agnd p2d p2d_b TGB
xi65 uin_n net082 avdd agnd p1d p1d_b TGB
xi64 vcm net082 avdd agnd p2d p2d_b TGB
xi60 vcm net0137 avdd agnd p2d p2d_b TGB
xi59 int1n net0137 avdd agnd p1d p1d_b TGB
xi13 amp_n opip avdd agnd p2 p2_b TGB
xi9 vthn net0161 avdd agnd p2d p2d_b TGB
xsw1 int2p net0155 avdd agnd p1d p1d_b TGB
xi2 int2n net0161 avdd agnd p1d p1d_b TGB
xsw4 vthp net0155 avdd agnd p2d p2d_b TGB
c20 opin net088 5e-15
cint1p_1 opin net0107 5e-15
cint1p_2 opin net0107 5e-15
c21 opip net082 5e-15
cint1n_1 opip net0137 5e-15
cint1n_2 opip net0137 5e-15
cintn opip net0161 5e-15
cintp opin net0155 5e-15
.ends adder_cmp_1b_CIFF2
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: int2_bhv
** View name: schematic
.subckt int2_bhv agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b inn inp iref outn outp pdn rst rst_b vcm vrefn vrefp
xop agnd avdd opin opip iref outn outp pdn vcm vcm fdopb
xi24 opin outp avdd agnd rst rst_b TGB
xi66 vcm net69 avdd agnd p2d p2d_b TGB
xsw5 inn net69 avdd agnd p1d p1d_b TGB
xi65 vcm net99 avdd agnd p2d p2d_b TGB
xsw6 inn_1 opip avdd agnd p2 p2_b TGB
xi25 opip outn avdd agnd rst rst_b TGB
xsw2 inp_1 opin avdd agnd p2 p2_b TGB
xsw3 vcm inp_1 avdd agnd p1 p1_b TGB
xsw1 inp net99 avdd agnd p1d p1d_b TGB
xsw7 vcm inn_1 avdd agnd p1 p1_b TGB
cfbp opin outp 10e-15
cfbn opip outn 10e-15
csn0 inn_1 net69 10e-15
csp0 inp_1 net99 10e-15
.ends int2_bhv
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: TOP_IADC_1b_bhv
** View name: schematic
xint1 agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b adcinn adcinp iref_1 int1n int1p pdn pvrefn pvrefn_b pvrefp pvrefp_b rst rst_b vcm vrefn vrefp int1_1b_bhv
xclk_fb agnd avdd dout p2d pvrefn pvrefn_b pvrefp pvrefp_b clk_fb_1bit
xquantizer_1b agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b dout iref_3 pdn adcinn adcinp vcm vcm vcm int1n int1p int2n int2p adder_cmp_1b_CIFF2
xint2 agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b int1n int1p iref_2 int2n int2p pdn rst rst_b vcm vrefn vrefp int2_bhv
*.END
