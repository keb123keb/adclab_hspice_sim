** Generated for: hspiceD
** Generated on: Sep 24 11:00:05 2019
** Design library name: ADC_SAR_DS_v1_zoom_adc_ych
** Design cell name: ADC_SAR_8bit_V4_4_DS_mod2lev5_ff
** Design view name: schematic


*****  .TEMP 25
*****  .OPTION
*****  +    ARTIST=2
*****  +    INGOLD=2
*****  +    MEASOUT=1
*****  +    PARHIER=LOCAL
*****  +    PSF=2

** Library name: cell_bhv
** Cell name: PMOS_B
** View name: schematic
*****  .subckt PMOS_B b d g s
*****  .ends PMOS_B
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: NMOS_B
** View name: schematic
*****  .subckt NMOS_B b d g s
*****  .ends NMOS_B
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: inv_bhv
** View name: schematic
.subckt inv_bhv dgnd vdd y yn
r1 net23 yn 10
c1 yn dgnd 5e-15
xp1 vdd net23 y vdd PMOS_B
xn1 dgnd net23 y dgnd NMOS_B
.ends inv_bhv
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: nand2_bhv
** View name: schematic
.subckt nand2_bhv dgnd vdd y1 y2 yn
xn1 dgnd yn y2 net8 NMOS_B
xi9 dgnd net8 y1 dgnd NMOS_B
xp1 vdd yn y1 vdd PMOS_B
xi10 vdd yn y2 vdd PMOS_B
.ends nand2_bhv
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: TGB
** View name: schematic
*****  .subckt TGB bi1 bi2 pwra sub t tn
*****  .ends TGB
** End of subcircuit definition.

** Library name: SAR_ADC_ych
** Cell name: DAC_SW
** View name: schematic
.subckt DAC_SW agnd avdd d dac d_b psamp psamp_b vin vrefn vrefp
xi7 agnd avdd pvrefn pvrefn_b inv_bhv
xi3 agnd avdd pvrefp pvrefp_b inv_bhv
xi20 agnd avdd net054 pvrefp inv_bhv
xi1 agnd avdd net049 pvrefn inv_bhv
xi2 agnd avdd psamp_b d_b net049 nand2_bhv
xi19 agnd avdd psamp_b d net054 nand2_bhv
xswp vrefp dac avdd agnd pvrefp pvrefp_b TGB
xswn vrefn dac avdd agnd pvrefn pvrefn_b TGB
xswin vin dac avdd agnd psamp psamp_b TGB
.ends DAC_SW
** End of subcircuit definition.

** Library name: SAR_ADC_ych
** Cell name: SA_DAC_8bit
** View name: schematic
.subckt SA_DAC_8bit agnd avdd d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 dac00 dac_0 dac_1 dac_2 dac_3 dac_4 dac_5 dac_6 dac_7 db_0 db_1 db_2 db_3 db_4 db_5 db_6 db_7 pdac psamp psamp_b vdac00 vin vrefn vrefp
xswdac_0 agnd avdd d_0 dac_0 db_0 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_1 agnd avdd d_1 dac_1 db_1 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_2 agnd avdd d_2 dac_2 db_2 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_3 agnd avdd d_3 dac_3 db_3 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_4 agnd avdd d_4 dac_4 db_4 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_5 agnd avdd d_5 dac_5 db_5 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_6 agnd avdd d_6 dac_6 db_6 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_7 agnd avdd d_7 dac_7 db_7 psamp psamp_b vin vrefn vrefp DAC_SW
xi1 agnd avdd pdac pdac_b inv_bhv
xswdac00 vdac00 dac00 avdd agnd pdac pdac_b TGB
xswvin vin dac00 avdd agnd psamp psamp_b TGB
.ends SA_DAC_8bit
** End of subcircuit definition.

** Library name: SAR_ADC_ych
** Cell name: SA_8bit_C_Array_with_DAC_monotonic_v4_unit_cap_two_stage
** View name: schematic
.subckt SA_8bit_C_Array_with_DAC_monotonic_v4_unit_cap_two_stage agnd avdd d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 db_0 db_1 db_2 db_3 db_4 db_5 db_6 db_7 pdac psamp psamp_b to_cmp vin vrefn vrefp
xsa_dac agnd avdd d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 net30 dac_0 dac_1 dac_2 dac_3 dac_4 dac_5 dac_6 dac_7 db_0 db_1 db_2 db_3 db_4 db_5 db_6 db_7 pdac psamp psamp_b net023 vrefp vrefn vrefp SA_DAC_8bit
xswvcmp vin to_cmp agnd avdd psamp psamp_b TGB
c8 to_cmp net038 12e-15
c0 net038 dac_0 12e-15
c2 net038 dac_2 24e-15
c1 net038 dac_1 12e-15
c3 net038 dac_3 48e-15
c4 net038 dac_4 96e-15
c7 to_cmp dac_7 48e-15
c5 to_cmp dac_5 12e-15
c6 to_cmp dac_6 24e-15
.ends SA_8bit_C_Array_with_DAC_monotonic_v4_unit_cap_two_stage
** End of subcircuit definition.

** Library name: SAR_ADC_ych
** Cell name: VCVS_CMP
** View name: schematic
*****  .subckt VCVS_CMP vm vout vp
*****  .ends VCVS_CMP
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: nor2_bhv
** View name: schematic
.subckt nor2_bhv dgnd vdd y1 y2 yn
xn1 dgnd yn y1 dgnd NMOS_B
xi9 dgnd yn y2 dgnd NMOS_B
xp1 vdd yn y2 net16 PMOS_B
xi10 vdd net16 y1 vdd PMOS_B
.ends nor2_bhv
** End of subcircuit definition.

** Library name: SAR_bhv
** Cell name: DFF_SET_RST
** View name: schematic
.subckt DFF_SET_RST q d clk dvdd dgnd set q_b rst
xi1 dgnd dvdd clk clkb inv_bhv
xi40 d dff1 dvdd dgnd clkb clk TGB
xi34 dff3 q_b dvdd dgnd clkb clk TGB
xi41 dff2 dff3 dvdd dgnd clk clkb TGB
xsw1 dff1 net41 dvdd dgnd clk clkb TGB
r1 net69 dff2 2
r0 net54 q 2
c3 q_b dgnd 100e-15
c2 net41 dgnd 100e-15
c4 q dgnd 100e-15
c1 dff2 dgnd 100e-15
xi42 dgnd dvdd dff2 rst net41 nor2_bhv
xi43 dgnd dvdd q set q_b nor2_bhv
xi31 dgnd dvdd dff1 set net69 nor2_bhv
xi37 dgnd dvdd dff3 rst net54 nor2_bhv
.ends DFF_SET_RST
** End of subcircuit definition.

** Library name: SAR_ADC_ych
** Cell name: SA_LOGIC_8bit_monotonic
** View name: schematic
.subckt SA_LOGIC_8bit_monotonic clk data_in d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 db_0 db_1 db_2 db_3 db_4 db_5 db_6 db_7 dgnd dvdd n_sw_0 n_sw_1 n_sw_2 n_sw_3 n_sw_4 n_sw_5 n_sw_6 n_sw_7 n_sw_b_0 n_sw_b_1 n_sw_b_2 n_sw_b_3 n_sw_b_4 n_sw_b_5 n_sw_b_6 n_sw_b_7 rst
xi36 dgnd dvdd data_in net383 inv_bhv
xi19 dgnd dvdd db_7 q7 n_sw_b_7 nor2_bhv
xi23 dgnd dvdd db_5 q5 n_sw_b_5 nor2_bhv
xi22 dgnd dvdd db_6 q6 n_sw_b_6 nor2_bhv
xi26 dgnd dvdd db_4 q4 n_sw_b_4 nor2_bhv
xi27 dgnd dvdd db_3 q3 n_sw_b_3 nor2_bhv
xi29 dgnd dvdd db_2 q2 n_sw_b_2 nor2_bhv
xi32 dgnd dvdd db_1 q1 n_sw_b_1 nor2_bhv
xi33 dgnd dvdd db_0 q0 n_sw_b_0 nor2_bhv
xi24 dgnd dvdd qb5 d_5 n_sw_5 nand2_bhv
xi20 dgnd dvdd d_7 qb7 n_sw_7 nand2_bhv
xi21 dgnd dvdd d_6 qb6 n_sw_6 nand2_bhv
xi25 dgnd dvdd qb4 d_4 n_sw_4 nand2_bhv
xi28 dgnd dvdd qb3 d_3 n_sw_3 nand2_bhv
xi30 dgnd dvdd qb2 d_2 n_sw_2 nand2_bhv
xi31 dgnd dvdd qb1 d_1 n_sw_1 nand2_bhv
xi34 dgnd dvdd qb0 d_0 n_sw_0 nand2_bhv
xdata3 d_3 net383 qb3 dvdd dgnd rst db_3 dgnd DFF_SET_RST
xdata2 d_2 net383 qb2 dvdd dgnd rst db_2 dgnd DFF_SET_RST
xdata1 d_1 net383 qb1 dvdd dgnd rst db_1 dgnd DFF_SET_RST
xdata0 d_0 net383 qb0 dvdd dgnd rst db_0 dgnd DFF_SET_RST
xdata5 d_5 net383 qb5 dvdd dgnd rst db_5 dgnd DFF_SET_RST
xrsh0 q0 q1 clk dvdd dgnd rst qb0 dgnd DFF_SET_RST
xrsh3 q3 q4 clk dvdd dgnd rst qb3 dgnd DFF_SET_RST
xrsh2 q2 q3 clk dvdd dgnd rst qb2 dgnd DFF_SET_RST
xrsh1 q1 q2 clk dvdd dgnd rst qb1 dgnd DFF_SET_RST
xrsh4 q4 q5 clk dvdd dgnd rst qb4 dgnd DFF_SET_RST
xdata7 d_7 net383 qb7 dvdd dgnd rst db_7 dgnd DFF_SET_RST
xrsh5 q5 q6 clk dvdd dgnd rst qb5 dgnd DFF_SET_RST
xdata6 d_6 net383 qb6 dvdd dgnd rst db_6 dgnd DFF_SET_RST
xdata4 d_4 net383 qb4 dvdd dgnd rst db_4 dgnd DFF_SET_RST
xrsh6 q6 q7 clk dvdd dgnd rst qb6 dgnd DFF_SET_RST
xrsh7 q7 dgnd clk dvdd dgnd rst qb7 dgnd DFF_SET_RST
.ends SA_LOGIC_8bit_monotonic
** End of subcircuit definition.

** Library name: SAR_ADC_ych
** Cell name: DFF_SET_RST
** View name: schematic
.subckt DFF_SET_RST_schematic q d clk dvdd dgnd set q_b rst
xi1 dgnd dvdd clk clkb inv_bhv
xi40 d dff1 dvdd dgnd clkb clk TGB
xi34 dff3 q_b dvdd dgnd clkb clk TGB
xi41 dff2 dff3 dvdd dgnd clk clkb TGB
xsw1 dff1 net41 dvdd dgnd clk clkb TGB
r1 net69 dff2 2
r0 net54 q 2
c3 q_b dgnd 100e-15
c2 net41 dgnd 100e-15
c4 q dgnd 100e-15
c1 dff2 dgnd 100e-15
xi42 dgnd dvdd dff2 rst net41 nor2_bhv
xi43 dgnd dvdd q set q_b nor2_bhv
xi31 dgnd dvdd dff1 set net69 nor2_bhv
xi37 dgnd dvdd dff3 rst net54 nor2_bhv
.ends DFF_SET_RST_schematic
** End of subcircuit definition.

** Library name: SAR_ADC_ych
** Cell name: ADC_SAR_diff_8bit_v4_monotonic_v4_unit_cap_two_stage
** View name: schematic
.subckt ADC_SAR_diff_8bit_v4_monotonic_v4_unit_cap_two_stage agnd avdd clk d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 dgnd dvdd psamp sa_7 sa_6 sa_5 sa_4 sa_3 sa_2 sa_1 sa_0 sa_b_7 sa_b_6 sa_b_5 sa_b_4 sa_b_3 sa_b_2 sa_b_1 sa_b_0 vinn vinp vrefn vrefp
xc_array_p agnd avdd db_0 db_1 db_2 db_3 db_4 db_5 db_6 db_7 d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 pdac psamp psamp_b cmp_inp vinp vrefn vrefp SA_8bit_C_Array_with_DAC_monotonic_v4_unit_cap_two_stage
xc_array_n agnd avdd n_sw_0 n_sw_1 n_sw_2 n_sw_3 n_sw_4 n_sw_5 n_sw_6 n_sw_7 n_sw_b_0 n_sw_b_1 n_sw_b_2 n_sw_b_3 n_sw_b_4 n_sw_b_5 n_sw_b_6 n_sw_b_7 pdac psamp psamp_b cmp_inn vinn vrefn vrefp SA_8bit_C_Array_with_DAC_monotonic_v4_unit_cap_two_stage
xcmp cmp_inn cmp_out cmp_inp VCVS_CMP
xsa_logic clk_b cmp_out db_0 db_1 db_2 db_3 db_4 db_5 db_6 db_7 d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 dgnd dvdd n_sw_0 n_sw_1 n_sw_2 n_sw_3 n_sw_4 n_sw_5 n_sw_6 n_sw_7 n_sw_b_0 n_sw_b_1 n_sw_b_2 n_sw_b_3 n_sw_b_4 n_sw_b_5 n_sw_b_6 n_sw_b_7 psamp SA_LOGIC_8bit_monotonic
xdffout_7 sa_7 d_7 psamp dvdd dgnd dgnd sa_b_7 dgnd DFF_SET_RST_schematic
xdffout_6 sa_6 d_6 psamp dvdd dgnd dgnd sa_b_6 dgnd DFF_SET_RST_schematic
xdffout_5 sa_5 d_5 psamp dvdd dgnd dgnd sa_b_5 dgnd DFF_SET_RST_schematic
xdffout_4 sa_4 d_4 psamp dvdd dgnd dgnd sa_b_4 dgnd DFF_SET_RST_schematic
xdffout_3 sa_3 d_3 psamp dvdd dgnd dgnd sa_b_3 dgnd DFF_SET_RST_schematic
xdffout_2 sa_2 d_2 psamp dvdd dgnd dgnd sa_b_2 dgnd DFF_SET_RST_schematic
xdffout_1 sa_1 d_1 psamp dvdd dgnd dgnd sa_b_1 dgnd DFF_SET_RST_schematic
xdffout_0 sa_0 d_0 psamp dvdd dgnd dgnd sa_b_0 dgnd DFF_SET_RST_schematic
xi7 dgnd dvdd psamp_b clk net23 nand2_bhv
xi28 dgnd dvdd clk clk_b inv_bhv
xi6 dgnd dvdd net23 pdac inv_bhv
xi5 dgnd dvdd psamp psamp_b inv_bhv
.ends ADC_SAR_diff_8bit_v4_monotonic_v4_unit_cap_two_stage
** End of subcircuit definition.

** Library name: adc_mod2_lev5_ff
** Cell name: Carray_8bit_sar_in
** View name: schematic
.subckt Carray_8bit_sar_in sar_cin_0 sar_cin_1 sar_cin_2 sar_cin_3 sar_cin_4 sar_cin_5 sar_cin_6 sar_cin_7 sar_dac_0 sar_dac_1 sar_dac_2 sar_dac_3 sar_dac_4 sar_dac_5 sar_dac_6 sar_dac_7
c_sar_n_1 sar_cin_1 sar_dac_1 312.5e-18
c_sar_n_2 sar_cin_2 sar_dac_2 625e-18
c_sar_n_7 sar_cin_7 sar_dac_7 20e-15
c_sar_n_6 sar_cin_6 sar_dac_6 10e-15
c_sar_n_5 sar_cin_5 sar_dac_5 5e-15
c_sar_n_4 sar_cin_4 sar_dac_4 2.5e-15
c_sar_n_0 sar_cin_0 sar_dac_0 156.25e-18
c_sar_n_3 sar_cin_3 sar_dac_3 1.25e-15
.ends Carray_8bit_sar_in
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: dac_int_1bit
** View name: schematic
.subckt dac_int_1bit agnd avdd dacn dacp pvrefn pvrefn_b pvrefp pvrefp_b vrefn vrefp
xi6 vrefn dacn avdd agnd pvrefp pvrefp_b TGB
xi7 vrefp dacn avdd agnd pvrefn pvrefn_b TGB
xi40 vrefp dacp avdd agnd pvrefp pvrefp_b TGB
xi41 vrefn dacp avdd agnd pvrefn pvrefn_b TGB
.ends dac_int_1bit
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: fdopb
** View name: schematic
*****  .subckt fdopb agnd avdd inn inp ir on op pdn vcm vcmfb
*****  .ends fdopb
** End of subcircuit definition.

** Library name: adc_mod2_lev5_ff
** Cell name: int1_with_lev5_dac_v2_8bit_sar_in
** View name: schematic
.subckt int1_with_lev5_dac_v2_8bit_sar_in agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b inn inp iref outn outp pdn pvrefn_0 pvrefn_1 pvrefn_2 pvrefn_3 pvrefn_b_0 pvrefn_b_1 pvrefn_b_2 pvrefn_b_3 pvrefp_0 pvrefp_1 pvrefp_2 pvrefp_3 pvrefp_b_0 pvrefp_b_1 pvrefp_b_2 pvrefp_b_3 rst rst_b sar_inn_0 sar_inn_1 sar_inn_2 sar_inn_3 sar_inn_4 sar_inn_5 sar_inn_6 sar_inn_7 sar_inp_0 sar_inp_1 sar_inp_2 sar_inp_3 sar_inp_4 sar_inp_5 sar_inp_6 sar_inp_7 vcm vrefn vrefp
xcarrayp sar_cinp_0 sar_cinp_1 sar_cinp_2 sar_cinp_3 sar_cinp_4 sar_cinp_5 sar_cinp_6 sar_cinp_7 sar_dacp_0 sar_dacp_1 sar_dacp_2 sar_dacp_3 sar_dacp_4 sar_dacp_5 sar_dacp_6 sar_dacp_7 Carray_8bit_sar_in
xcarrayn sar_cinn_0 sar_cinn_1 sar_cinn_2 sar_cinn_3 sar_cinn_4 sar_cinn_5 sar_cinn_6 sar_cinn_7 sar_dacn_0 sar_dacn_1 sar_dacn_2 sar_dacn_3 sar_dacn_4 sar_dacn_5 sar_dacn_6 sar_dacn_7 Carray_8bit_sar_in
xdac_0 agnd avdd dacn_0 dacp_0 pvrefn_0 pvrefn_b_0 pvrefp_0 pvrefp_b_0 vrefn vrefp dac_int_1bit
xdac_1 agnd avdd dacn_1 dacp_1 pvrefn_1 pvrefn_b_1 pvrefp_1 pvrefp_b_1 vrefn vrefp dac_int_1bit
xdac_2 agnd avdd dacn_2 dacp_2 pvrefn_2 pvrefn_b_2 pvrefp_2 pvrefp_b_2 vrefn vrefp dac_int_1bit
xdac_3 agnd avdd dacn_3 dacp_3 pvrefn_3 pvrefn_b_3 pvrefp_3 pvrefp_b_3 vrefn vrefp dac_int_1bit
cfbp_0 opip outp 10e-15
cfbp_1 opip outp 10e-15
cfbp_2 opip outp 10e-15
cfbp_3 opip outp 10e-15
c1_0 cinp dacp_0 10e-15
c1_1 cinp dacp_1 10e-15
c1_2 cinp dacp_2 10e-15
c1_3 cinp dacp_3 10e-15
c2_0 cinn dacn_0 10e-15
c2_1 cinn dacn_1 10e-15
c2_2 cinn dacn_2 10e-15
c2_3 cinn dacn_3 10e-15
cfbn_0 opin outn 10e-15
cfbn_1 opin outn 10e-15
cfbn_2 opin outn 10e-15
cfbn_3 opin outn 10e-15
xsw3 vcm cinp avdd agnd p1 p1_b TGB
xsw7 vcm cinn avdd agnd p1 p1_b TGB
xsw4_0 sar_cinp_0 opip avdd agnd p2 p2_b TGB
xsw4_1 sar_cinp_1 opip avdd agnd p2 p2_b TGB
xsw4_2 sar_cinp_2 opip avdd agnd p2 p2_b TGB
xsw4_3 sar_cinp_3 opip avdd agnd p2 p2_b TGB
xsw4_4 sar_cinp_4 opip avdd agnd p2 p2_b TGB
xsw4_5 sar_cinp_5 opip avdd agnd p2 p2_b TGB
xsw4_6 sar_cinp_6 opip avdd agnd p2 p2_b TGB
xsw4_7 sar_cinp_7 opip avdd agnd p2 p2_b TGB
xsw_sar_inp_0 sar_inp_0 sar_dacp_0 avdd agnd p2d p2d_b TGB
xsw_sar_inp_1 sar_inp_1 sar_dacp_1 avdd agnd p2d p2d_b TGB
xsw_sar_inp_2 sar_inp_2 sar_dacp_2 avdd agnd p2d p2d_b TGB
xsw_sar_inp_3 sar_inp_3 sar_dacp_3 avdd agnd p2d p2d_b TGB
xsw_sar_inp_4 sar_inp_4 sar_dacp_4 avdd agnd p2d p2d_b TGB
xsw_sar_inp_5 sar_inp_5 sar_dacp_5 avdd agnd p2d p2d_b TGB
xsw_sar_inp_6 sar_inp_6 sar_dacp_6 avdd agnd p2d p2d_b TGB
xsw_sar_inp_7 sar_inp_7 sar_dacp_7 avdd agnd p2d p2d_b TGB
xsw_sar_inn_0 sar_inn_0 sar_dacn_0 avdd agnd p2d p2d_b TGB
xsw_sar_inn_1 sar_inn_1 sar_dacn_1 avdd agnd p2d p2d_b TGB
xsw_sar_inn_2 sar_inn_2 sar_dacn_2 avdd agnd p2d p2d_b TGB
xsw_sar_inn_3 sar_inn_3 sar_dacn_3 avdd agnd p2d p2d_b TGB
xsw_sar_inn_4 sar_inn_4 sar_dacn_4 avdd agnd p2d p2d_b TGB
xsw_sar_inn_5 sar_inn_5 sar_dacn_5 avdd agnd p2d p2d_b TGB
xsw_sar_inn_6 sar_inn_6 sar_dacn_6 avdd agnd p2d p2d_b TGB
xsw_sar_inn_7 sar_inn_7 sar_dacn_7 avdd agnd p2d p2d_b TGB
xswinn_0 inn dacn_0 avdd agnd p1d p1d_b TGB
xswinn_1 inn dacn_1 avdd agnd p1d p1d_b TGB
xswinn_2 inn dacn_2 avdd agnd p1d p1d_b TGB
xswinn_3 inn dacn_3 avdd agnd p1d p1d_b TGB
xsw5_0 sar_cinn_0 opin avdd agnd p2 p2_b TGB
xsw5_1 sar_cinn_1 opin avdd agnd p2 p2_b TGB
xsw5_2 sar_cinn_2 opin avdd agnd p2 p2_b TGB
xsw5_3 sar_cinn_3 opin avdd agnd p2 p2_b TGB
xsw5_4 sar_cinn_4 opin avdd agnd p2 p2_b TGB
xsw5_5 sar_cinn_5 opin avdd agnd p2 p2_b TGB
xsw5_6 sar_cinn_6 opin avdd agnd p2 p2_b TGB
xsw5_7 sar_cinn_7 opin avdd agnd p2 p2_b TGB
xsw2 cinp opip avdd agnd p2 p2_b TGB
xsw6 cinn opin avdd agnd p2 p2_b TGB
xi12 outn opin avdd agnd rst rst_b TGB
xi13 outp opip avdd agnd rst rst_b TGB
xswinp_0 inp dacp_0 avdd agnd p1d p1d_b TGB
xswinp_1 inp dacp_1 avdd agnd p1d p1d_b TGB
xswinp_2 inp dacp_2 avdd agnd p1d p1d_b TGB
xswinp_3 inp dacp_3 avdd agnd p1d p1d_b TGB
xop agnd avdd opip opin iref outn outp pdn vcm vcm fdopb
.ends int1_with_lev5_dac_v2_8bit_sar_in
** End of subcircuit definition.

** Library name: adc_mod2_lev5_ff
** Cell name: int2
** View name: schematic
.subckt int2 agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b inn inp iref outn outp pdn rst rst_b vcm
c0 cinp dacp 10e-15
c3 cinn dacn 10e-15
c4 opip outp 10e-15
c5 opin outn 10e-15
xi65 vcm dacp avdd agnd p2d p2d_b TGB
xsw7 vcm cinn avdd agnd p1 p1_b TGB
xsw3 vcm cinp avdd agnd p1 p1_b TGB
xswinn_0 inn dacn avdd agnd p1d p1d_b TGB
xswinn_1 inn dacn avdd agnd p1d p1d_b TGB
xswinn_2 inn dacn avdd agnd p1d p1d_b TGB
xswinn_3 inn dacn avdd agnd p1d p1d_b TGB
xswinp_0 inp dacp avdd agnd p1d p1d_b TGB
xswinp_1 inp dacp avdd agnd p1d p1d_b TGB
xswinp_2 inp dacp avdd agnd p1d p1d_b TGB
xswinp_3 inp dacp avdd agnd p1d p1d_b TGB
xsw2 cinp opip avdd agnd p2 p2_b TGB
xsw6 cinn opin avdd agnd p2 p2_b TGB
xi6 outn opin avdd agnd rst rst_b TGB
xi9 outp opip avdd agnd rst rst_b TGB
xi66 vcm dacn avdd agnd p2d p2d_b TGB
xop agnd avdd opip opin iref outn outp pdn vcm vcm fdopb
.ends int2
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: preamp_cmp_b
** View name: schematic
*****  .subckt preamp_cmp_b agnd avdd inn inp ir on op pdn vcm vcmfb
*****  .ends preamp_cmp_b
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: Dlatch
** View name: schematic
.subckt Dlatch q d clk clkb dvdd dgnd
xi2 dgnd dvdd net017 q inv_bhv
xi1 dgnd dvdd net22 net8 inv_bhv
c0 q dgnd 5e-15
c1 net017 dgnd 5e-15
r1 net8 net017 2
xi29 d net22 dvdd dgnd clk clkb TGB
xsw1 net22 q dvdd dgnd clkb clk TGB
.ends Dlatch
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: dff
** View name: schematic
.subckt dff q d clk clkb dvdd dgnd
xi13 net275 d clkb clk dvdd dgnd Dlatch
xi14 q net275 clk clkb dvdd dgnd Dlatch
.ends dff
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: amp_cmp
** View name: schematic
*****  .subckt amp_cmp vm vout vp
*****  .ends amp_cmp
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: cmp_clk
** View name: schematic
.subckt cmp_clk agnd avdd clk clk_b inn inp y
xdff y net22 clk clk_b avdd agnd dff
xpreamp inn net22 inp amp_cmp
.ends cmp_clk
** End of subcircuit definition.

** Library name: adc_mod2_lev5_ff
** Cell name: adder_cmp_1b_CIFF2
** View name: schematic
.subckt adder_cmp_1b_CIFF2 agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b d iref pdn uin_n uin_p vcm vthn vthp int1n int1p int2n int2p
xpreamp_bhv agnd avdd opin opip iref amp_n amp_p pdn vcm vcm preamp_cmp_b
xcmp3 agnd avdd p1_b p1 amp_n amp_p d_b cmp_clk
xi1 agnd avdd d_b d inv_bhv
xi52 amp_p opin avdd agnd p2 p2_b TGB
xi63 vcm net088 avdd agnd p2d p2d_b TGB
xi62 uin_p net088 avdd agnd p1d p1d_b TGB
xi55 int1p net0107 avdd agnd p1d p1d_b TGB
xi56 vcm net0107 avdd agnd p2d p2d_b TGB
xi65 uin_n net082 avdd agnd p1d p1d_b TGB
xi64 vcm net082 avdd agnd p2d p2d_b TGB
xi60 vcm net0137 avdd agnd p2d p2d_b TGB
xi59 int1n net0137 avdd agnd p1d p1d_b TGB
xi13 amp_n opip avdd agnd p2 p2_b TGB
xi9 vthn net0161 avdd agnd p2d p2d_b TGB
xsw1 int2p net0155 avdd agnd p1d p1d_b TGB
xi2 int2n net0161 avdd agnd p1d p1d_b TGB
xsw4 vthp net0155 avdd agnd p2d p2d_b TGB
c20 opin net088 10e-15
cint1p_1 opin net0107 10e-15
cint1p_2 opin net0107 10e-15
c21 opip net082 10e-15
cint1n_1 opip net0137 10e-15
cint1n_2 opip net0137 10e-15
cintn opip net0161 10e-15
cintp opin net0155 10e-15
.ends adder_cmp_1b_CIFF2
** End of subcircuit definition.

** Library name: adc_mod2_lev5_ff
** Cell name: vth_5Lev
** View name: schematic
.subckt vth_5Lev vrefn vrefp vthp_0 vthp_1 vthp_2 vthp_3
r25 vthp_2 vthp_3 50e3
r9 vrefn vthp_0 50e3
r18 vrefp vthp_3 50e3
r8 vrefn vthp_0 50e3
r3 vthp_1 vthp_2 50e3
r2 vthp_0 vthp_1 50e3
r1 vrefp vthp_3 50e3
.ends vth_5Lev
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: clk_fb_1bit
** View name: schematic
.subckt clk_fb_1bit agnd avdd d p2 pvrefn pvrefn_b pvrefp pvrefp_b
xi64 agnd avdd pvrefn pvrefn_b inv_bhv
xi20 agnd avdd net43 pvrefp inv_bhv
xi60 agnd avdd net48 pvrefn inv_bhv
xi59 agnd avdd d d_b inv_bhv
xi63 agnd avdd pvrefp pvrefp_b inv_bhv
xi62 agnd avdd p2 d_b net48 nand2_bhv
xi19 agnd avdd p2 d net43 nand2_bhv
.ends clk_fb_1bit
** End of subcircuit definition.

** Library name: adc_mod2_lev5_ff
** Cell name: adc_mod2_lev5_ff_v2_8bit_sar_in
** View name: schematic
.subckt adc_mod2_lev5_ff_v2_8bit_sar_in agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b dgnd dout_0 dout_1 dout_2 dout_3 dvdd inn inp iref_1 iref_2 iref_cmp_0 iref_cmp_1 iref_cmp_2 iref_cmp_3 out_int2_n out_int2_p pdn rst rst_b sar_inn_0 sar_inn_1 sar_inn_2 sar_inn_3 sar_inn_4 sar_inn_5 sar_inn_6 sar_inn_7 sar_inp_0 sar_inp_1 sar_inp_2 sar_inp_3 sar_inp_4 sar_inp_5 sar_inp_6 sar_inp_7 vcm vrefn vrefp
xint1 agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b inn inp iref_1 out_int1_n out_int1_p pdn pvrefn_0 pvrefn_1 pvrefn_2 pvrefn_3 pvrefn_b_0 pvrefn_b_1 pvrefn_b_2 pvrefn_b_3 pvrefp_0 pvrefp_1 pvrefp_2 pvrefp_3 pvrefp_b_0 pvrefp_b_1 pvrefp_b_2 pvrefp_b_3 rst rst_b sar_inn_0 sar_inn_1 sar_inn_2 sar_inn_3 sar_inn_4 sar_inn_5 sar_inn_6 sar_inn_7 sar_inp_0 sar_inp_1 sar_inp_2 sar_inp_3 sar_inp_4 sar_inp_5 sar_inp_6 sar_inp_7 vcm vrefn vrefp int1_with_lev5_dac_v2_8bit_sar_in
xint2 agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b out_int1_n out_int1_p iref_2 out_int2_n out_int2_p pdn rst rst_b vcm int2
xquantizer_1b_0 agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b dout_0 iref_cmp_0 pdn inn inp vcm vthp_3 vthp_0 out_int1_n out_int1_p out_int2_n out_int2_p adder_cmp_1b_CIFF2
xquantizer_1b_1 agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b dout_1 iref_cmp_1 pdn inn inp vcm vthp_2 vthp_1 out_int1_n out_int1_p out_int2_n out_int2_p adder_cmp_1b_CIFF2
xquantizer_1b_2 agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b dout_2 iref_cmp_2 pdn inn inp vcm vthp_1 vthp_2 out_int1_n out_int1_p out_int2_n out_int2_p adder_cmp_1b_CIFF2
xquantizer_1b_3 agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b dout_3 iref_cmp_3 pdn inn inp vcm vthp_0 vthp_3 out_int1_n out_int1_p out_int2_n out_int2_p adder_cmp_1b_CIFF2
xvth vrefn vrefp vthp_0 vthp_1 vthp_2 vthp_3 vth_5Lev
xclk_fb_0 agnd avdd dout_0 p2d pvrefn_0 pvrefn_b_0 pvrefp_0 pvrefp_b_0 clk_fb_1bit
xclk_fb_1 agnd avdd dout_1 p2d pvrefn_1 pvrefn_b_1 pvrefp_1 pvrefp_b_1 clk_fb_1bit
xclk_fb_2 agnd avdd dout_2 p2d pvrefn_2 pvrefn_b_2 pvrefp_2 pvrefp_b_2 clk_fb_1bit
xclk_fb_3 agnd avdd dout_3 p2d pvrefn_3 pvrefn_b_3 pvrefp_3 pvrefp_b_3 clk_fb_1bit
.ends adc_mod2_lev5_ff_v2_8bit_sar_in
** End of subcircuit definition.

** Library name: ADC_SAR_DS_v1_zoom_adc_ych
** Cell name: ADC_SAR_8bit_V4_4_DS_mod2lev5_ff
** View name: schematic
xsar agnd avdd clk_sar d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 dgnd dvdd psamp sa_7 sa_6 sa_5 sa_4 sa_3 sa_2 sa_1 sa_0 sa_b_7 sa_b_6 sa_b_5 sa_b_4 sa_b_3 sa_b_2 sa_b_1 sa_b_0 inn inp vrefn vrefp ADC_SAR_diff_8bit_v4_monotonic_v4_unit_cap_two_stage
xds agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b dgnd dsout_0 dsout_1 dsout_2 dsout_3 dvdd inn inp iref_1 iref_2 iref_cmp_0 iref_cmp_1 iref_cmp_2 iref_cmp_3 out_int2_n out_int2_p pdn rst rst_b sa_b_0 sa_b_1 sa_b_2 sa_b_3 sa_b_4 sa_b_5 sa_b_6 sa_b_7 sa_0 sa_1 sa_2 sa_3 sa_4 sa_5 sa_6 sa_7 vcm vrefn vrefp adc_mod2_lev5_ff_v2_8bit_sar_in
*****  .END
