** Generated for: hspiceD
** Generated on: May  7 11:24:11 2019
** Design library name: myfirstlib
** Design cell name: 1int_1bit_fb
** Design view name: schematic


.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    MEASOUT=1
+    PARHIER=LOCAL
+    PSF=2

** Library name: cell_bhv
** Cell name: PMOS_B
** View name: schematic
.subckt PMOS_B b d g s
.ends PMOS_B
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: NMOS_B
** View name: schematic
.subckt NMOS_B b d g s
.ends NMOS_B
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: inv_bhv
** View name: schematic
.subckt inv_bhv dgnd vdd y yn
r1 net23 yn 10
c1 yn dgnd 5e-15
xp1 vdd net23 y vdd PMOS_B
xn1 dgnd net23 y dgnd NMOS_B
.ends inv_bhv
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: TGB
** View name: schematic
.subckt TGB bi1 bi2 pwra sub t tn
.ends TGB
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: Dlatch
** View name: schematic
.subckt Dlatch q d clk clkb dvdd dgnd
xi2 dgnd dvdd net017 q inv_bhv
xi1 dgnd dvdd net22 net8 inv_bhv
c0 q dgnd 5e-15
c1 net017 dgnd 5e-15
r1 net8 net017 2
xi29 d net22 dvdd dgnd clk clkb TGB
xsw1 net22 q dvdd dgnd clkb clk TGB
.ends Dlatch
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: dff
** View name: schematic
.subckt dff q d clk clkb dvdd dgnd
xi13 net275 d clkb clk dvdd dgnd Dlatch
xi14 q net275 clk clkb dvdd dgnd Dlatch
.ends dff
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: amp_cmp
** View name: schematic
.subckt amp_cmp vm vout vp
.ends amp_cmp
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: cmp_clk
** View name: schematic
.subckt cmp_clk agnd avdd clk clk_b inn inp y
xdff y net22 clk clk_b avdd agnd dff
xpreamp inn net22 inp amp_cmp
.ends cmp_clk
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: preamp_cmp_b
** View name: schematic
.subckt preamp_cmp_b agnd avdd inn inp ir on op pdn vcm vcmfb
.ends preamp_cmp_b
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: nand2_bhv
** View name: schematic
.subckt nand2_bhv dgnd vdd y1 y2 yn
xn1 dgnd yn y2 net8 NMOS_B
xi9 dgnd net8 y1 dgnd NMOS_B
xp1 vdd yn y1 vdd PMOS_B
xi10 vdd yn y2 vdd PMOS_B
.ends nand2_bhv
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: clk_fb_1bit
** View name: schematic
.subckt clk_fb_1bit agnd avdd d p2 pvrefn pvrefn_b pvrefp pvrefp_b
xi64 agnd avdd pvrefn pvrefn_b inv_bhv
xi20 agnd avdd net43 pvrefp inv_bhv
xi60 agnd avdd net48 pvrefn inv_bhv
xi59 agnd avdd d d_b inv_bhv
xi63 agnd avdd pvrefp pvrefp_b inv_bhv
xi62 agnd avdd p2 d_b net48 nand2_bhv
xi19 agnd avdd p2 d net43 nand2_bhv
.ends clk_fb_1bit
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: dac_int_1bit
** View name: schematic
.subckt dac_int_1bit agnd avdd dacn dacp pvrefn pvrefn_b pvrefp pvrefp_b vrefn vrefp
xi6 vrefn dacn avdd agnd pvrefp pvrefp_b TGB
xi7 vrefp dacn avdd agnd pvrefn pvrefn_b TGB
xi40 vrefp dacp avdd agnd pvrefp pvrefp_b TGB
xi41 vrefn dacp avdd agnd pvrefn pvrefn_b TGB
.ends dac_int_1bit
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: fdopb
** View name: schematic
.subckt fdopb agnd avdd inn inp ir on op pdn vcm vcmfb
.ends fdopb
** End of subcircuit definition.

** Library name: myfirstlib
** Cell name: 1int_1bit_fb
** View name: schematic
cintn opin_cmp acn_cmp 5e-15
cintp opip_cmp acp_cmp 5e-15
xi14 agnd avdd d_b dout inv_bhv
xcmp3 agnd avdd p1_b p1 amp_n amp_p d_b cmp_clk
xpreamp_bhv agnd avdd opip_cmp opin_cmp iref_2 amp_n amp_p pdn vcm vcm preamp_cmp_b
xclk_fb agnd avdd dout p2d pvrefn pvrefn_b pvrefp pvrefp_b clk_fb_1bit
xi10 agnd avdd dacn dacp pvrefn pvrefn_b pvrefp pvrefp_b vrefn vrefp dac_int_1bit
xi8 agnd avdd opip opin iref_1 out_int1_n out_int1_p pdn vcm vcm fdopb
xi9 vthn acn_cmp avdd agnd p2d p2d_b TGB
xi16 out_int1_n acn_cmp avdd agnd p1d p1d_b TGB
xi0 inp dacp avdd agnd p1d p1d_b TGB
xi1 dacn inn avdd agnd p1d p1d_b TGB
xi2 opin cinn avdd agnd p2 p2_b TGB
xi3 cinp opip avdd agnd p2 p2_b TGB
xi5 vcm cinn avdd agnd p1 p1_b TGB
xi7 vcm cinp avdd agnd p1 p1_b TGB
xi13 out_int1_p opip avdd agnd rst rst_b TGB
xi12 out_int1_n opin avdd agnd rst rst_b TGB
xsw4 vthp acp_cmp avdd agnd p2d p2d_b TGB
xsw1 out_int1_p acp_cmp avdd agnd p1d p1d_b TGB
xi52 amp_p opip_cmp avdd agnd p2 p2_b TGB
xi15 amp_n opin_cmp avdd agnd p2 p2_b TGB
cfbn_1 opin out_int1_n 100e-15
cfbn_2 opin out_int1_n 100e-15
cfbn_3 opin out_int1_n 100e-15
c2 cinn dacn 100e-15
c1 cinp dacp 100e-15
cfbp_1 opip out_int1_p 100e-15
cfbp_2 opip out_int1_p 100e-15
cfbp_3 opip out_int1_p 100e-15
.END
