** Generated for: hspiceD
** Generated on: Jan 11 04:42:23 2020
** Design library name: ADC_DS_SAR_v1_extented_range_ych
** Design cell name: ADC_DS_mod2bit1_ff_SAR_10bit_v2_split_c
** Design view name: schematic
*****  .PARAM k kp


*****  .TEMP 25
*****  .OPTION
*****  +    ARTIST=2
*****  +    INGOLD=2
*****  +    MEASOUT=1
*****  +    PARHIER=LOCAL
*****  +    PSF=2

** Library name: cell_bhv
** Cell name: PMOS_B
** View name: schematic
*****  .subckt PMOS_B b d g s
*****  .ends PMOS_B
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: NMOS_B
** View name: schematic
*****  .subckt NMOS_B b d g s
*****  .ends NMOS_B
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: inv_bhv
** View name: schematic
.subckt inv_bhv dgnd vdd y yn
r1 net23 yn 10
c1 yn dgnd 5e-15
xp1 vdd net23 y vdd PMOS_B
xn1 dgnd net23 y dgnd NMOS_B
.ends inv_bhv
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: TGB
** View name: schematic
*****  .subckt TGB bi1 bi2 pwra sub t tn
*****  .ends TGB
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: nor2_bhv
** View name: schematic
.subckt nor2_bhv dgnd vdd y1 y2 yn
xn1 dgnd yn y1 dgnd NMOS_B
xi9 dgnd yn y2 dgnd NMOS_B
xp1 vdd yn y2 net16 PMOS_B
xi10 vdd net16 y1 vdd PMOS_B
.ends nor2_bhv
** End of subcircuit definition.

** Library name: SAR_bhv
** Cell name: DFF_SET_RST
** View name: schematic
.subckt DFF_SET_RST q d clk dvdd dgnd set q_b rst
xi1 dgnd dvdd clk clkb inv_bhv
xi40 d dff1 dvdd dgnd clkb clk TGB
xi34 dff3 q_b dvdd dgnd clkb clk TGB
xi41 dff2 dff3 dvdd dgnd clk clkb TGB
xsw1 dff1 net41 dvdd dgnd clk clkb TGB
r1 net69 dff2 2
r0 net54 q 2
c3 q_b dgnd 100e-15
c2 net41 dgnd 100e-15
c4 q dgnd 100e-15
c1 dff2 dgnd 100e-15
xi42 dgnd dvdd dff2 rst net41 nor2_bhv
xi43 dgnd dvdd q set q_b nor2_bhv
xi31 dgnd dvdd dff1 set net69 nor2_bhv
xi37 dgnd dvdd dff3 rst net54 nor2_bhv
.ends DFF_SET_RST
** End of subcircuit definition.

** Library name: SAR_ADC_ych
** Cell name: SA_LOGIC_10bit
** View name: schematic
.subckt SA_LOGIC_10bit clk comp d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 d_8 d_9 db_0 db_1 db_2 db_3 db_4 db_5 db_6 db_7 db_8 db_9 dgnd dvdd rst
xdata9 d_9 comp d_8 dvdd dgnd q9 db_9 dgnd DFF_SET_RST
xdata8 d_8 comp d_7 dvdd dgnd q8 db_8 rst DFF_SET_RST
xrsh8 q8 q9 clk dvdd dgnd dgnd net086 rst DFF_SET_RST
xrsh9 q9 dgnd clk dvdd dgnd rst net078 dgnd DFF_SET_RST
xrsh00 q00 q0 clk dvdd dgnd dgnd net0150 rst DFF_SET_RST
xdata3 d_3 comp d_2 dvdd dgnd q3 db_3 rst DFF_SET_RST
xdata2 d_2 comp d_1 dvdd dgnd q2 db_2 rst DFF_SET_RST
xdata1 d_1 comp d_0 dvdd dgnd q1 db_1 rst DFF_SET_RST
xdata00 net089 dgnd dgnd dvdd dgnd q00 net060 rst DFF_SET_RST
xdata0 d_0 comp net089 dvdd dgnd q0 db_0 rst DFF_SET_RST
xdata5 d_5 comp d_4 dvdd dgnd q5 db_5 rst DFF_SET_RST
xrsh0 q0 q1 clk dvdd dgnd dgnd net0158 rst DFF_SET_RST
xrsh3 q3 q4 clk dvdd dgnd dgnd net0166 rst DFF_SET_RST
xrsh2 q2 q3 clk dvdd dgnd dgnd net0174 rst DFF_SET_RST
xrsh1 q1 q2 clk dvdd dgnd dgnd net0182 rst DFF_SET_RST
xrsh4 q4 q5 clk dvdd dgnd dgnd net0190 rst DFF_SET_RST
xdata7 d_7 comp d_6 dvdd dgnd q7 db_7 rst DFF_SET_RST
xrsh5 q5 q6 clk dvdd dgnd dgnd net0198 rst DFF_SET_RST
xdata6 d_6 comp d_5 dvdd dgnd q6 db_6 rst DFF_SET_RST
xdata4 d_4 comp d_3 dvdd dgnd q4 db_4 rst DFF_SET_RST
xrsh6 q6 q7 clk dvdd dgnd dgnd net0206 rst DFF_SET_RST
xrsh7 q7 q8 clk dvdd dgnd dgnd net0214 rst DFF_SET_RST
.ends SA_LOGIC_10bit
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: nand2_bhv
** View name: schematic
.subckt nand2_bhv dgnd vdd y1 y2 yn
xn1 dgnd yn y2 net8 NMOS_B
xi9 dgnd net8 y1 dgnd NMOS_B
xp1 vdd yn y1 vdd PMOS_B
xi10 vdd yn y2 vdd PMOS_B
.ends nand2_bhv
** End of subcircuit definition.

** Library name: SAR_ADC_ych
** Cell name: DAC_SW
** View name: schematic
.subckt DAC_SW agnd avdd d dac d_b psamp psamp_b vin vrefn vrefp
xi7 agnd avdd pvrefn pvrefn_b inv_bhv
xi3 agnd avdd pvrefp pvrefp_b inv_bhv
xi20 agnd avdd net054 pvrefp inv_bhv
xi1 agnd avdd net049 pvrefn inv_bhv
xi2 agnd avdd psamp_b d_b net049 nand2_bhv
xi19 agnd avdd psamp_b d net054 nand2_bhv
xswp vrefp dac avdd agnd pvrefp pvrefp_b TGB
xswn vrefn dac avdd agnd pvrefn pvrefn_b TGB
xswin vin dac avdd agnd psamp psamp_b TGB
.ends DAC_SW
** End of subcircuit definition.

** Library name: SAR_ADC_ych
** Cell name: SA_DAC_10bit
** View name: schematic
.subckt SA_DAC_10bit agnd avdd d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 dac00 dac_0 dac_1 dac_2 dac_3 dac_4 dac_5 dac_6 dac_7 db_0 db_1 db_2 db_3 db_4 db_5 db_6 db_7 pdac psamp psamp_b vdac00 vin vrefn vrefp d_8 d_9 dac_8 dac_9 db_8 db_9
xswdac_0 agnd avdd d_0 dac_0 db_0 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_1 agnd avdd d_1 dac_1 db_1 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_2 agnd avdd d_2 dac_2 db_2 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_3 agnd avdd d_3 dac_3 db_3 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_4 agnd avdd d_4 dac_4 db_4 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_5 agnd avdd d_5 dac_5 db_5 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_6 agnd avdd d_6 dac_6 db_6 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_7 agnd avdd d_7 dac_7 db_7 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_8 agnd avdd d_8 dac_8 db_8 psamp psamp_b vin vrefn vrefp DAC_SW
xswdac_9 agnd avdd d_9 dac_9 db_9 psamp psamp_b vin vrefn vrefp DAC_SW
xi1 agnd avdd pdac pdac_b inv_bhv
xswdac00 vdac00 dac00 avdd agnd pdac pdac_b TGB
xswvin vin dac00 avdd agnd psamp psamp_b TGB
.ends SA_DAC_10bit
** End of subcircuit definition.

** Library name: SAR_ADC_ych
** Cell name: SA_10bit_C_Array_with_DAC_two_stage
** View name: schematic
.subckt SA_10bit_C_Array_with_DAC_two_stage agnd avdd d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 db_0 db_1 db_2 db_3 db_4 db_5 db_6 db_7 pdac psamp psamp_b to_cmp vcm vdac00 vinp vrefn vrefp d_8 d_9 db_8 db_9
xsa_dac agnd avdd d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 dac00 dac_0 dac_1 dac_2 dac_3 dac_4 dac_5 dac_6 dac_7 db_0 db_1 db_2 db_3 db_4 db_5 db_6 db_7 pdac psamp psamp_b vdac00 vinp vrefn vrefp d_8 d_9 dac_8 dac_9 db_8 db_9 SA_DAC_10bit
xi2 vcm to_cmp agnd avdd psamp psamp_b TGB
cp1 vrefp net47 '(12e-15/k)*kp'
cp2 vrefp to_cmp '(12e-15/k)*kp'
c00 net47 dac00 '12e-15/k'
c9 to_cmp dac_9 '192e-15/k'
c4 net47 dac_4 '192e-15/k'
**c0 to_cmp net47 '12.387096774194e-15/k'
c0 to_cmp net47 '12e-15/k'
c1 net47 dac_0 '12e-15/k'
c2 net47 dac_2 '48e-15/k'
c3 net47 dac_1 '24e-15/k'
c5 net47 dac_3 '96e-15/k'
c6 to_cmp dac_5 '12e-15/k'
c8 to_cmp dac_8 '96e-15/k'
c7 to_cmp dac_6 '24e-15/k'
c10 to_cmp dac_7 '48e-15/k'
.ends SA_10bit_C_Array_with_DAC_two_stage
** End of subcircuit definition.

** Library name: SAR_ADC_ych
** Cell name: VCVS_CMP
** View name: schematic
*****  .subckt VCVS_CMP vm vout vp
*****  .ends VCVS_CMP
** End of subcircuit definition.

** Library name: SAR_ADC_ych
** Cell name: DFF_SET_RST
** View name: schematic
.subckt DFF_SET_RST_schematic q d clk dvdd dgnd set q_b rst
xi1 dgnd dvdd clk clkb inv_bhv
xi40 d dff1 dvdd dgnd clkb clk TGB
xi34 dff3 q_b dvdd dgnd clkb clk TGB
xi41 dff2 dff3 dvdd dgnd clk clkb TGB
xsw1 dff1 net41 dvdd dgnd clk clkb TGB
r1 net69 dff2 2
r0 net54 q 2
c3 q_b dgnd 100e-15
c2 net41 dgnd 100e-15
c4 q dgnd 100e-15
c1 dff2 dgnd 100e-15
xi42 dgnd dvdd dff2 rst net41 nor2_bhv
xi43 dgnd dvdd q set q_b nor2_bhv
xi31 dgnd dvdd dff1 set net69 nor2_bhv
xi37 dgnd dvdd dff3 rst net54 nor2_bhv
.ends DFF_SET_RST_schematic
** End of subcircuit definition.

** Library name: cell_bhv
** Cell name: Dlatch
** View name: schematic
.subckt Dlatch q d clk clkb dvdd dgnd
xi2 dgnd dvdd net017 q inv_bhv
xi1 dgnd dvdd net22 net8 inv_bhv
c0 q dgnd 5e-15
c1 net017 dgnd 5e-15
r1 net8 net017 2
xi29 d net22 dvdd dgnd clk clkb TGB
xsw1 net22 q dvdd dgnd clkb clk TGB
.ends Dlatch
** End of subcircuit definition.

** Library name: SAR_ADC_ych
** Cell name: ADC_SAR_diff_10bit_v2_two_stage
** View name: schematic
.subckt ADC_SAR_diff_10bit_v2_two_stage agnd avdd clk d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 d_8 d_9 dgnd dvdd psamp sa_9 sa_8 sa_7 sa_6 sa_5 sa_4 sa_3 sa_2 sa_1 sa_0 sa_b_9 sa_b_8 sa_b_7 sa_b_6 sa_b_5 sa_b_4 sa_b_3 sa_b_2 sa_b_1 sa_b_0 vinn vinp vrefn vrefp
xi27 pdac_b cmp_out d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 d_8 d_9 db_0 db_1 db_2 db_3 db_4 db_5 db_6 db_7 db_8 db_9 dgnd dvdd psamp SA_LOGIC_10bit
xc_array_p agnd avdd d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 db_0 db_1 db_2 db_3 db_4 db_5 db_6 db_7 pdac psamp psamp_b cmp_inn vcm vrefn vinp vrefn vrefp d_8 d_9 db_8 db_9 SA_10bit_C_Array_with_DAC_two_stage
xc_array_n agnd avdd d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 db_0 db_1 db_2 db_3 db_4 db_5 db_6 db_7 pdac psamp psamp_b cmp_inp vcm vrefp vinn vrefp vrefn d_8 d_9 db_8 db_9 SA_10bit_C_Array_with_DAC_two_stage
xi24 cmp_inn cmp_diff cmp_inp VCVS_CMP
xdffout_9 sa_9 d_9 psamp dvdd dgnd dgnd sa_b_9 dgnd DFF_SET_RST_schematic
xdffout_8 sa_8 d_8 psamp dvdd dgnd dgnd sa_b_8 dgnd DFF_SET_RST_schematic
xdffout_7 sa_7 d_7 psamp dvdd dgnd dgnd sa_b_7 dgnd DFF_SET_RST_schematic
xdffout_6 sa_6 d_6 psamp dvdd dgnd dgnd sa_b_6 dgnd DFF_SET_RST_schematic
xdffout_5 sa_5 d_5 psamp dvdd dgnd dgnd sa_b_5 dgnd DFF_SET_RST_schematic
xdffout_4 sa_4 d_4 psamp dvdd dgnd dgnd sa_b_4 dgnd DFF_SET_RST_schematic
xdffout_3 sa_3 d_3 psamp dvdd dgnd dgnd sa_b_3 dgnd DFF_SET_RST_schematic
xdffout_2 sa_2 d_2 psamp dvdd dgnd dgnd sa_b_2 dgnd DFF_SET_RST_schematic
xdffout_1 sa_1 d_1 psamp dvdd dgnd dgnd sa_b_1 dgnd DFF_SET_RST_schematic
xdffout_0 sa_0 d_0 psamp dvdd dgnd dgnd sa_b_0 dgnd DFF_SET_RST_schematic
xi7 dgnd dvdd psamp_b clk net69 nand2_bhv
xi8 dgnd dvdd pdac pdac_b inv_bhv
xi6 dgnd dvdd net69 pdac inv_bhv
xi5 dgnd dvdd psamp psamp_b inv_bhv
xcmplatch cmp_out cmp_diff pdac pdac_b dvdd dgnd Dlatch
.ends ADC_SAR_diff_10bit_v2_two_stage
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: dac_int_1bit
** View name: schematic
.subckt dac_int_1bit agnd avdd dacn dacp pvrefn pvrefn_b pvrefp pvrefp_b vrefn vrefp
xi6 vrefn dacn avdd agnd pvrefp pvrefp_b TGB
xi7 vrefp dacn avdd agnd pvrefn pvrefn_b TGB
xi40 vrefp dacp avdd agnd pvrefp pvrefp_b TGB
xi41 vrefn dacp avdd agnd pvrefn pvrefn_b TGB
.ends dac_int_1bit
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: fdopb
** View name: schematic
*****  .subckt fdopb agnd avdd inn inp ir on op pdn vcm vcmfb
*****  .ends fdopb
** End of subcircuit definition.

** Library name: adc_mod2_bit1_ff
** Cell name: int1_G103_with_1b_dac
** View name: schematic
.subckt int1_G103_with_1b_dac agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b inn inp iref outn outp pdn pvrefn pvrefn_b pvrefp pvrefp_b rst rst_b vcm vrefn vrefp
xdac agnd avdd dacn dacp pvrefn pvrefn_b pvrefp pvrefp_b vrefn vrefp dac_int_1bit
cfbp_1 opip outp 10e-15
cfbp_2 opip outp 10e-15
cfbp_3 opip outp 10e-15
c1 cinp dacp 10e-15
c2 cinn dacn 10e-15
cfbn_1 opin outn 10e-15
cfbn_2 opin outn 10e-15
cfbn_3 opin outn 10e-15
xsw3 vcm cinp avdd agnd p1 p1_b TGB
xsw7 vcm cinn avdd agnd p1 p1_b TGB
xswinn inn dacn avdd agnd p1d p1d_b TGB
xsw2 cinp opip avdd agnd p2 p2_b TGB
xsw6 cinn opin avdd agnd p2 p2_b TGB
xi12 outn opin avdd agnd rst rst_b TGB
xi13 outp opip avdd agnd rst rst_b TGB
xswinp inp dacp avdd agnd p1d p1d_b TGB
xop agnd avdd opip opin iref outn outp pdn vcm vcm fdopb
.ends int1_G103_with_1b_dac
** End of subcircuit definition.

** Library name: adc_mod2_bit1_ff
** Cell name: int2
** View name: schematic
.subckt int2 agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b inn inp iref outn outp pdn rst rst_b vcm
c0 cinp dacp 10e-15
c3 cinn dacn 10e-15
cfbp opip outp 10e-15
cfbn opin outn 10e-15
xi65 vcm dacp avdd agnd p2d p2d_b TGB
xsw7 vcm cinn avdd agnd p1 p1_b TGB
xsw3 vcm cinp avdd agnd p1 p1_b TGB
xswinn inn dacn avdd agnd p1d p1d_b TGB
xswinp inp dacp avdd agnd p1d p1d_b TGB
xsw2 cinp opip avdd agnd p2 p2_b TGB
xsw6 cinn opin avdd agnd p2 p2_b TGB
xi6 outn opin avdd agnd rst rst_b TGB
xi9 outp opip avdd agnd rst rst_b TGB
xi66 vcm dacn avdd agnd p2d p2d_b TGB
xop agnd avdd opip opin iref outn outp pdn vcm vcm fdopb
.ends int2
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: preamp_cmp_b
** View name: schematic
*****  .subckt preamp_cmp_b agnd avdd inn inp ir on op pdn vcm vcmfb
*****  .ends preamp_cmp_b
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: dff
** View name: schematic
.subckt dff q d clk clkb dvdd dgnd
xi13 net275 d clkb clk dvdd dgnd Dlatch
xi14 q net275 clk clkb dvdd dgnd Dlatch
.ends dff
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: amp_cmp
** View name: schematic
*****  .subckt amp_cmp vm vout vp
*****  .ends amp_cmp
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: cmp_clk
** View name: schematic
.subckt cmp_clk agnd avdd clk clk_b inn inp y
xdff y net22 clk clk_b avdd agnd dff
xpreamp inn net22 inp amp_cmp
.ends cmp_clk
** End of subcircuit definition.

** Library name: adc_mod2_bit1_ff
** Cell name: adder_cmp_1b_CIFF2
** View name: schematic
.subckt adder_cmp_1b_CIFF2 agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b d iref pdn uin_n uin_p vcm vthn vthp int1n int1p int2n int2p
xpreamp_bhv agnd avdd opin opip iref amp_n amp_p pdn vcm vcm preamp_cmp_b
xcmp3 agnd avdd p1_b p1 amp_n amp_p d_b cmp_clk
xi1 agnd avdd d_b d inv_bhv
xi52 amp_p opin avdd agnd p2 p2_b TGB
xi63 vcm net088 avdd agnd p2d p2d_b TGB
xi62 uin_p net088 avdd agnd p1d p1d_b TGB
xi55 int1p net0107 avdd agnd p1d p1d_b TGB
xi56 vcm net0107 avdd agnd p2d p2d_b TGB
xi65 uin_n net082 avdd agnd p1d p1d_b TGB
xi64 vcm net082 avdd agnd p2d p2d_b TGB
xi60 vcm net0137 avdd agnd p2d p2d_b TGB
xi59 int1n net0137 avdd agnd p1d p1d_b TGB
xi13 amp_n opip avdd agnd p2 p2_b TGB
xi9 vthn net0161 avdd agnd p2d p2d_b TGB
xsw1 int2p net0155 avdd agnd p1d p1d_b TGB
xi2 int2n net0161 avdd agnd p1d p1d_b TGB
xsw4 vthp net0155 avdd agnd p2d p2d_b TGB
c20 opin net088 10e-15
cint1p_1 opin net0107 10e-15
cint1p_2 opin net0107 10e-15
cint1p_3 opin net0107 10e-15
cint1p_4 opin net0107 10e-15
cint1p_5 opin net0107 10e-15
cint1p_6 opin net0107 10e-15
c21 opip net082 10e-15
cint1n_1 opip net0137 10e-15
cint1n_2 opip net0137 10e-15
cint1n_3 opip net0137 10e-15
cint1n_4 opip net0137 10e-15
cint1n_5 opip net0137 10e-15
cint1n_6 opip net0137 10e-15
cintn_1 opip net0161 10e-15
cintn_2 opip net0161 10e-15
cintn_3 opip net0161 10e-15
cintp_1 opin net0155 10e-15
cintp_2 opin net0155 10e-15
cintp_3 opin net0155 10e-15
.ends adder_cmp_1b_CIFF2
** End of subcircuit definition.

** Library name: ET710_ADC_bhv
** Cell name: clk_fb_1bit
** View name: schematic
.subckt clk_fb_1bit agnd avdd d p2 pvrefn pvrefn_b pvrefp pvrefp_b
xi64 agnd avdd pvrefn pvrefn_b inv_bhv
xi20 agnd avdd net43 pvrefp inv_bhv
xi60 agnd avdd net48 pvrefn inv_bhv
xi59 agnd avdd d d_b inv_bhv
xi63 agnd avdd pvrefp pvrefp_b inv_bhv
xi62 agnd avdd p2 d_b net48 nand2_bhv
xi19 agnd avdd p2 d net43 nand2_bhv
.ends clk_fb_1bit
** End of subcircuit definition.

** Library name: adc_mod2_bit1_ff
** Cell name: adc_mod2_bit1_ff
** View name: schematic
.subckt adc_mod2_bit1_ff agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b dgnd dout dvdd inn inp iref_1 iref_2 iref_3 out_int2_n out_int2_p pdn rst rst_b vcm vrefn vrefp
xint1 agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b inn inp iref_1 out_int1_n out_int1_p pdn pvrefn pvrefn_b pvrefp pvrefp_b rst rst_b vcm vrefn vrefp int1_G103_with_1b_dac
xint2 agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b out_int1_n out_int1_p iref_2 out_int2_n out_int2_p pdn rst rst_b vcm int2
xquantizer agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b dout iref_3 pdn inn inp vcm vcm vcm out_int1_n out_int1_p out_int2_n out_int2_p adder_cmp_1b_CIFF2
xclk_fb agnd avdd dout p2d pvrefn pvrefn_b pvrefp pvrefp_b clk_fb_1bit
.ends adc_mod2_bit1_ff
** End of subcircuit definition.

** Library name: ADC_DS_SAR_v1_extented_range_ych
** Cell name: ADC_DS_mod2bit1_ff_SAR_10bit_v2_split_c
** View name: schematic
xsar agnd avdd clk_sar d_0 d_1 d_2 d_3 d_4 d_5 d_6 d_7 d_8 d_9 dgnd dvdd psamp sa_9 sa_8 sa_7 sa_6 sa_5 sa_4 sa_3 sa_2 sa_1 sa_0 sa_b_9 sa_b_8 sa_b_7 sa_b_6 sa_b_5 sa_b_4 sa_b_3 sa_b_2 sa_b_1 sa_b_0 residualxg1o3_n residualxg1o3_p vrefn vrefp ADC_SAR_diff_10bit_v2_two_stage
xds agnd avdd p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b dgnd ds_out dvdd inn inp iref_1 iref_2 iref_3 residualxg1o3_n residualxg1o3_p pdn rst rst_b vcm vrefn vrefp adc_mod2_bit1_ff
*****  .END
